--- This file will include: Receiver, Transmitter, BaudRateGenerator ---