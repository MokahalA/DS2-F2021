--- This file will include: UART FSM ---